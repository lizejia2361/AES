module Sub_Bytes(
    input wire [127:0] state, // 128位输入状态
    output wire [127:0] subbed_state // 128位输出状态，经过S盒字节代换后的结果
);

// S盒定义
function [7:0] S;
    input [7:0] x;
    begin
        case (x)
            8'd0  : S = 8'h63;
            8'd1  : S = 8'h7c;
            8'd2  : S = 8'h77;
            8'd3  : S = 8'h7b;
            8'd4  : S = 8'hf2;
            8'd5  : S = 8'h6b;
            8'd6  : S = 8'h6f;
            8'd7  : S = 8'hc5;
            8'd8  : S = 8'h30;
            8'd9  : S = 8'h01;
            8'd10 : S = 8'h67;
            8'd11 : S = 8'h2b;
            8'd12 : S = 8'hfe;
            8'd13 : S = 8'hd7;
            8'd14 : S = 8'hab;
            8'd15 : S = 8'h76;
            8'd16 : S = 8'hca;
            8'd17 : S = 8'h82;
            8'd18 : S = 8'hc9;
            8'd19 : S = 8'h7d;
            8'd20 : S = 8'hfa;
            8'd21 : S = 8'h59;
            8'd22 : S = 8'h47;
            8'd23 : S = 8'hf0;
            8'd24 : S = 8'had;
            8'd25 : S = 8'hd4;
            8'd26 : S = 8'ha2;
            8'd27 : S = 8'haf;
            8'd28 : S = 8'h9c;
            8'd29 : S = 8'ha4;
            8'd30 : S = 8'h72;
            8'd31 : S = 8'hc0;
            8'd32 : S = 8'hb7;
            8'd33 : S = 8'hfd;
            8'd34 : S = 8'h93;
            8'd35 : S = 8'h26;
            8'd36 : S = 8'h36;
            8'd37 : S = 8'h3f;
            8'd38 : S = 8'hf7;
            8'd39 : S = 8'hcc;
            8'd40 : S = 8'h34;
            8'd41 : S = 8'ha5;
            8'd42 : S = 8'he5;
            8'd43 : S = 8'hf1;
            8'd44 : S = 8'h71;
            8'd45 : S = 8'hd8;
            8'd46 : S = 8'h31;
            8'd47 : S = 8'h15;
            8'd48 : S = 8'h04;
            8'd49 : S = 8'hc7;
            8'd50 : S = 8'h23;
            8'd51 : S = 8'hc3;
            8'd52 : S = 8'h18;
            8'd53 : S = 8'h96;
            8'd54 : S = 8'h05;
            8'd55 : S = 8'h9a;
            8'd56 : S = 8'h07;
            8'd57 : S = 8'h12;
            8'd58 : S = 8'h80;
            8'd59 : S = 8'he2;
            8'd60 : S = 8'heb;
            8'd61 : S = 8'h27;
            8'd62 : S = 8'hb2;
            8'd63 : S = 8'h75;
            8'd64 : S = 8'h09;
            8'd65 : S = 8'h83;
            8'd66 : S = 8'h2c;
            8'd67 : S = 8'h1a;
            8'd68 : S = 8'h1b;
            8'd69 : S = 8'h6e;
            8'd70 : S = 8'h5a;
            8'd71 : S = 8'ha0;
            8'd72 : S = 8'h52;
            8'd73 : S = 8'h3b;
            8'd74 : S = 8'hd6;
            8'd75 : S = 8'hb3;
            8'd76 : S = 8'h29;
            8'd77 : S = 8'he3;
            8'd78 : S = 8'h2f;
            8'd79 : S = 8'h84;
            8'd80 : S = 8'h53;
            8'd81 : S = 8'hd1;
            8'd82 : S = 8'h00;
            8'd83 : S = 8'hed;
            8'd84 : S = 8'h20;
            8'd85 : S = 8'hfc;
            8'd86 : S = 8'hb1;
            8'd87 : S = 8'h5b;
            8'd88 : S = 8'h6a;
            8'd89 : S = 8'hcb;
            8'd90 : S = 8'hbe;
            8'd91 : S = 8'h39;
            8'd92 : S = 8'h4a;
            8'd93 : S = 8'h4c;
            8'd94 : S = 8'h58;
            8'd95 : S = 8'hcf;
            8'd96 : S = 8'hd0;
            8'd97 : S = 8'hef;
            8'd98 : S = 8'haa;
            8'd99 : S = 8'hfb;
            8'd100: S = 8'h43;
            8'd101: S = 8'h4d;
            8'd102: S = 8'h33;
            8'd103: S = 8'h85;
            8'd104: S = 8'h45;
            8'd105: S = 8'hf9;
            8'd106: S = 8'h02;
            8'd107: S = 8'h7f;
            8'd108: S = 8'h50;
            8'd109: S = 8'h3c;
            8'd110: S = 8'h9f;
            8'd111: S = 8'ha8;
            8'd112: S = 8'h51;
            8'd113: S = 8'ha3;
            8'd114: S = 8'h40;
            8'd115: S = 8'h8f;
            8'd116: S = 8'h92;
            8'd117: S = 8'h9d;
            8'd118: S = 8'h38;
            8'd119: S = 8'hf5;
            8'd120: S = 8'hbc;
            8'd121: S = 8'hb6;
            8'd122: S = 8'hda;
            8'd123: S = 8'h21;
            8'd124: S = 8'h10;
            8'd125: S = 8'hff;
            8'd126: S = 8'hf3;
            8'd127: S = 8'hd2;
            8'd128: S = 8'hcd;
            8'd129: S = 8'h0c;
            8'd130: S = 8'h13;
            8'd131: S = 8'hec;
            8'd132: S = 8'h5f;
            8'd133: S = 8'h97;
            8'd134: S = 8'h44;
            8'd135: S = 8'h17;
            8'd136: S = 8'hc4;
            8'd137: S = 8'ha7;
            8'd138: S = 8'h7e;
            8'd139: S = 8'h3d;
            8'd140: S = 8'h64;
            8'd141: S = 8'h5d;
            8'd142: S = 8'h19;
            8'd143: S = 8'h73;
            8'd144: S = 8'h60;
            8'd145: S = 8'h81;
            8'd146: S = 8'h4f;
            8'd147: S = 8'hdc;
            8'd148: S = 8'h22;
            8'd149: S = 8'h2a;
            8'd150: S = 8'h90;
            8'd151: S = 8'h88;
            8'd152: S = 8'h46;
            8'd153: S = 8'hee;
            8'd154: S = 8'hb8;
            8'd155: S = 8'h14;
            8'd156: S = 8'hde;
            8'd157: S = 8'h5e;
            8'd158: S = 8'h0b;
            8'd159: S = 8'hdb;
            8'd160: S = 8'he0; 
            8'd161: S = 8'h32; 
            8'd162: S = 8'h3a; 
            8'd163: S = 8'h0a; 
            8'd164: S = 8'h49; 
            8'd165: S = 8'h06; 
            8'd166: S = 8'h24; 
            8'd167: S = 8'h5c; 
            8'd168: S = 8'hc2; 
            8'd169: S = 8'hd3; 
            8'd170: S = 8'hac; 
            8'd171: S = 8'h62; 
            8'd172: S = 8'h91; 
            8'd173: S = 8'h95; 
            8'd174: S = 8'he4; 
            8'd175: S = 8'h79; 
            8'd176: S = 8'he7; 
            8'd177: S = 8'hc8; 
            8'd178: S = 8'h37; 
            8'd179: S = 8'h6d; 
            8'd180: S = 8'h8d; 
            8'd181: S = 8'hd5; 
            8'd182: S = 8'h4e; 
            8'd183: S = 8'ha9; 
            8'd184: S = 8'h6c; 
            8'd185: S = 8'h56; 
            8'd186: S = 8'hf4; 
            8'd187: S = 8'hea; 
            8'd188: S = 8'h65; 
            8'd189: S = 8'h7a; 
            8'd190: S = 8'hae; 
            8'd191: S = 8'h08; 
            8'd192: S = 8'hba; 
            8'd193: S = 8'h78; 
            8'd194: S = 8'h25; 
            8'd195: S = 8'h2e; 
            8'd196: S = 8'h1c; 
            8'd197: S = 8'ha6; 
            8'd198: S = 8'hb4; 
            8'd199: S = 8'hc6; 
            8'd200: S = 8'he8; 
            8'd201: S = 8'hdd; 
            8'd202: S = 8'h74; 
            8'd203: S = 8'h1f; 
            8'd204: S = 8'h4b; 
            8'd205: S = 8'hbd; 
            8'd206: S = 8'h8b; 
            8'd207: S = 8'h8a; 
            8'd208: S = 8'h70; 
            8'd209: S = 8'h3e; 
            8'd210: S = 8'hb5; 
            8'd211: S = 8'h66; 
            8'd212: S = 8'h48; 
            8'd213: S = 8'h03; 
            8'd214: S = 8'hf6; 
            8'd215: S = 8'h0e; 
            8'd216: S = 8'h61; 
            8'd217: S = 8'h35; 
            8'd218: S = 8'h57; 
            8'd219: S = 8'hb9; 
            8'd220: S = 8'h86; 
            8'd221: S = 8'hc1; 
            8'd222: S = 8'h1d; 
            8'd223: S = 8'h9e; 
            8'd224: S = 8'he1; 
            8'd225: S = 8'hf8; 
            8'd226: S = 8'h98; 
            8'd227: S = 8'h11; 
            8'd228: S = 8'h69; 
            8'd229: S = 8'hd9; 
            8'd230: S = 8'h8e; 
            8'd231: S = 8'h94; 
            8'd232: S = 8'h9b; 
            8'd233: S = 8'h1e; 
            8'd234: S = 8'h87; 
            8'd235: S = 8'he9; 
            8'd236: S = 8'hce; 
            8'd237: S = 8'h55; 
            8'd238: S = 8'h28; 
            8'd239: S = 8'hdf; 
            8'd240: S = 8'h8c; 
            8'd241: S = 8'ha1;
            8'd242: S = 8'h89; 
            8'd243: S = 8'h0d; 
            8'd244: S = 8'hbf; 
            8'd245: S = 8'he6; 
            8'd246: S = 8'h42; 
            8'd247: S = 8'h68;
            8'd248: S = 8'h41; 
            8'd249: S = 8'h99; 
            8'd250: S = 8'h2d; 
            8'd251: S = 8'h0f; 
            8'd252: S = 8'hb0; 
            8'd253: S = 8'h54;
            8'd254: S = 8'hbb;
            8'd255: S = 8'd16;
            default: S = 8'd0;
        endcase
    end
endfunction

// 将128位输入状态分解为16个8位字节，并分别进行S盒代换
wire [7:0] byte0, byte1, byte2, byte3, byte4, byte5, byte6, byte7,
           byte8, byte9, byte10, byte11, byte12, byte13, byte14, byte15;

assign byte0 = state[7:0];
assign byte1 = state[15:8];
assign byte2 = state[23:16];
assign byte3 = state[31:24];
assign byte4 = state[39:32];
assign byte5 = state[47:40];
assign byte6 = state[55:48];
assign byte7 = state[63:56];
assign byte8 = state[71:64];
assign byte9 = state[79:72];
assign byte10 = state[87:80];
assign byte11 = state[95:88];
assign byte12 = state[103:96];
assign byte13 = state[111:104];
assign byte14 = state[119:112];
assign byte15 = state[127:120];

// 应用S盒代换
wire [7:0] subbed_byte0, subbed_byte1, subbed_byte2, subbed_byte3,
           subbed_byte4, subbed_byte5, subbed_byte6, subbed_byte7,
           subbed_byte8, subbed_byte9, subbed_byte10, subbed_byte11,
           subbed_byte12, subbed_byte13, subbed_byte14, subbed_byte15;

assign subbed_byte0 = S(byte0);
assign subbed_byte1 = S(byte1);
assign subbed_byte2 = S(byte2);
assign subbed_byte3 = S(byte3);
assign subbed_byte4 = S(byte4);
assign subbed_byte5 = S(byte5);
assign subbed_byte6 = S(byte6);
assign subbed_byte7 = S(byte7);
assign subbed_byte8 = S(byte8);
assign subbed_byte9 = S(byte9);
assign subbed_byte10 = S(byte10);
assign subbed_byte11 = S(byte11);
assign subbed_byte12 = S(byte12);
assign subbed_byte13 = S(byte13);
assign subbed_byte14 = S(byte14);
assign subbed_byte15 = S(byte15);

// 将代换后的字节重新组合成128位输出状态
assign subbed_state = {subbed_byte15, subbed_byte14, subbed_byte13, subbed_byte12,
                       subbed_byte11, subbed_byte10, subbed_byte9, subbed_byte8,
                       subbed_byte7, subbed_byte6, subbed_byte5, subbed_byte4,
                       subbed_byte3, subbed_byte2, subbed_byte1, subbed_byte0};

endmodule